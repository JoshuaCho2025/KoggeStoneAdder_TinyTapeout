`default_nettype none
`timescale 1ns / 1ps

/* This testbench instantiates the 8-bit Kogge-Stone adder module 
   and provides convenient wires for driving and testing with cocotb.
*/
module tb ();

  // Dump the signals to a VCD file. You can view it with gtkwave.
  initial begin
    $dumpfile("tb.vcd");
    $dumpvars(0, tb);
    #1;
  end

  // Wire up the inputs and outputs:
  reg clk;
  reg rst_n;
  reg ena;
  reg [7:0] a, b;
  reg [7:0] uio_in;
  wire [7:0] sum;
  wire carry_out;
  wire [7:0] uio_out;
  wire [7:0] uio_oe;
`ifdef GL_TEST
  wire VPWR = 1'b1;
  wire VGND = 1'b0;
`endif

  // Instantiate the 8-bit Kogge-Stone adder module:
  tt_um_koggestone_adder8 user_project (

      // Include power ports for the Gate Level test:
`ifdef GL_TEST
      .VPWR(VPWR),
      .VGND(VGND),
`endif

      .ui_in  ({b, a}),          // 8-bit input (concatenated a and b)
      .uo_out (sum),             // 8-bit sum output
      .uio_in (uio_in),          // IOs: Input path
      .uio_out(uio_out),         // IOs: Output path
      .uio_oe (uio_oe),          // IOs: Enable path (active high: 0=input, 1=output)
      .ena    (ena),             // Enable - goes high when design is selected
      .clk    (clk),             // Clock
      .rst_n  (rst_n)            // Active-low reset
  );

endmodule
